library verilog;
use verilog.vl_types.all;
entity Problem_3_vlg_vec_tst is
end Problem_3_vlg_vec_tst;
