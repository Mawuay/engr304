library verilog;
use verilog.vl_types.all;
entity Problem8_vlg_vec_tst is
end Problem8_vlg_vec_tst;
