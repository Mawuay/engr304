library verilog;
use verilog.vl_types.all;
entity Problem4_vlg_vec_tst is
end Problem4_vlg_vec_tst;
