library verilog;
use verilog.vl_types.all;
entity ThunderBird_vlg_vec_tst is
end ThunderBird_vlg_vec_tst;
