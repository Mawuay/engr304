library verilog;
use verilog.vl_types.all;
entity Problem4 is
    port(
        f2              : out    vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        x4              : in     vl_logic;
        f1              : out    vl_logic
    );
end Problem4;
