library ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.fulladd_package.all ; -- declare package here
