library verilog;
use verilog.vl_types.all;
entity Problem_3 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        F               : out    vl_logic
    );
end Problem_3;
